`timescale 1ns/1ps

module full_adder (
    input a, b, cin,
    output sumo, cout
    );

    assign sumo = a ^ b ^ cin;
    assign cout = (a & b) | (b & cin) | (cin & a);
endmodule

module parallel_adder (
    input [3:0] A, B,
    input carry_in,
    output [3:0] sum,
    output carry
    );  

    wire [2:0] c;
    full_adder fa0 (A[0], B[0], carry_in, sum[0], c[0]);
    full_adder fa1 (A[1], B[1], c[0], sum[1], c[1]);            // aint this called instantiation?
    full_adder fa2 (A[2], B[2], c[1], sum[2], c[2]);
    full_adder fa3 (A[3], B[3], c[2], sum[3], carry);

endmodule       
